/////////////////////////////////////////////////////////////////////
// ---------------------- IVCAD 2020 Spring ---------------------- //
// ---------------------- Editor : Claire C ---------------------- //
// ---------------------- Version : v.1.00  ---------------------- //
// ---------------------- Date : 2020.02.05 ---------------------- //
// ----------------------        adder      ---------------------- //
/////////////////////////////////////////////////////////////////////

module sat_adder(in0, in1, in2, sum);

input  signed[33:0]	in0, in1, in2;
output signed[15:0]	sum;

wire signed[35:0]temp=(in0+in1+in2);
assign sum=($signed(temp)>$signed(36'd255))?16'd255:($signed(temp)<$signed(36'd0))?16'd0:temp[15:0];

endmodule
